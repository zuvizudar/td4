module rom(dout, addr);
	output [7:0] dout;
	input [3:0] addr;

	reg[7:0] mem[15:0];

	initial begin
		mem[4'b0000] <= 8'b1011_0111;
		mem[4'b0001] <= 8'b0000_0001;	
		mem[4'b0010] <= 8'b1110_0001;	
		mem[4'b0011] <= 8'b0000_0001;	
		mem[4'b0100] <= 8'b1110_0011;	
		mem[4'b0101] <= 8'b1011_0110;	
		mem[4'b0110] <= 8'b0000_0001;	
		mem[4'b0111] <= 8'b1110_0101;	
		mem[4'b1000] <= 8'b0000_0001;	
		mem[4'b1001] <= 8'b0000_1000;
		mem[4'b1010] <= 8'b1011_0100;
		mem[4'b1011] <= 8'b1001_0000;
		mem[4'b1100] <= 8'b0000_0001;
		mem[4'b1101] <= 8'b1110_1010;
		mem[4'b1110] <= 8'b1011_1000;
		mem[4'b1111] <= 8'b1111_1111;
	end

	assign dout = mem[addr];
endmodule